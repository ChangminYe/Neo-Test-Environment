// Parameters
`define CLKS_PER_BIT 868    // Num
`define GLOBAL_NEURON 2**16 // Num

